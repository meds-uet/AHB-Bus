// Parameters declaration

parameter DATA_WIDTH = 32;
parameter ADDR_WIDTH = 32;

parameter MASTER_NUM = 3;
