// Copyright 2025 Maktab-e-Digital Systems Lahore.
// Licensed under the Apache License, Version 2.0, see LICENSE file for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: 
// This module contains the parameters for AHB bus.
//
//
// Author: Muhammad Yousaf and Ali Tahir
// Date:   29-July-2025


parameter integer NUM_MASTERS = 4;
parameter integer NUM_SLAVES = 4;
parameter integer DATA_WIDTH = 32;
parameter integer ADDR_WIDTH = 32;